//A console for playing a fighting game
//The goal of the game is knocking out your opponent whit a variation of attacks
//interface: leds for feedback, reset button, VGA interface, switches for settings 

module console(iCLK_50, iKEY, iSW, oVGA_R, oVGA_G, oVGA_B, oVGA_HS, oVGA_VS, oVGA_CLOCK, oVGA_SYNC_N, oVGA_BLANK_N, oLEDR, GPIO_0);

//input and output values
	//clock, switches and buttons
	input iCLK_50;
	input [0:0] iKEY;
	input [17:0] iSW;
	input [4:0] GPIO_0;
	
	//VGA
	output  oVGA_CLOCK; 
	output [9:0] oVGA_R, oVGA_G, oVGA_B;
	output oVGA_HS, oVGA_VS;
	output oVGA_SYNC_N; 
	output oVGA_BLANK_N;
	output [17:0] oLEDR;
	
	//testing
	//wire test;
	assign oLEDR[9:0] = controller1;
	
	//define interfaces
	//reset button
	wire reset;
	assign reset = ~iKEY[0];

	//VGA with picture processing unit (ppsu)
	//attributes is used by the statemachine to ajust the moving sprites in the ppu
	//wire [] attributes;
	wire hsync, vsync;
	assign oVGA_CLOCK = clock;
	assign oVGA_SYNC_N = 1'b0;
	assign oVGA_HS = hsync; assign oVGA_VS = vsync;
	assign oVGA_BLANK_N = hsync & vsync;
	
	//connection between statemachine and ppu

	wire [9:0] red, green, blue;
	
	wire [63:0] sprites;
	wire [0:0] statics;
	
	ppu picture_proc_unit(.clock(clock), .reset(reset), .red(red), .green(green), .blue(blue), .hsync(hsync), .vsync(vsync), 
						  .sprites(sprites), .statics(statics), .test(iSW[1:0]));

	assign oVGA_R = red;
	assign oVGA_G = green;
	assign oVGA_B = blue;
	
	//the game statemachine
	wire [9:0] controller1;
	wire [9:0] controller2;
	statemachine sm(.clock(clock), .reset(reset), .controller1(controller1), .controller2(controller2), 
					.sprites(sprites), .statics(statics), .test(oLEDR[17]));
	
	//input
	ps2_connect inputcontroller(.clock(clock), .reset(reset), .GPIO_0(GPIO_0), .c1(controller1), .c2(controller2));
	
	//rom
	//not yet implemented
	
	//clock signal with pll - 108Mhz
	wire clock;
	pll pll(reset, iCLK_50, clock);


endmodule 