module statemachine(clock, reset, controls, sprites, statics, offset_x, offset_y, update);

input clock, reset;
input [17:0] controls;
input update;

output [179:0] sprites;
output [131:0] statics;
output [11:0] offset_x, offset_y;

assign sprites = 0;
assign statics = 0;
assign offset_x = 0;
assign offset_y = 0;

//declaration of the statemachine

endmodule 